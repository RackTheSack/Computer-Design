/*
  Eric Villasenor
  evillase@gmail.com

  register file test bench
*/

// mapped needs this
`include "register_file_if.vh"

// mapped timing needs this. 1ns is too fast
`timescale 1 ns / 1 ns

module register_file_tb;

  parameter PERIOD = 10;

  logic CLK = 0, nRST;

  // test vars
  int v1 = 1;
  int v2 = 4721;
  int v3 = 25119;

  // clock
  always #(PERIOD/2) CLK++;

  // interface
  register_file_if rfif ();
  // test program
  test #(.PERIOD (PERIOD)) PROG(
    CLK,
    nRST,
    rfif
  );
  // DUT
`ifndef MAPPED
  register_file DUT(CLK, nRST, rfif);
`else
  register_file DUT(
    .\rfif.rdat2 (rfif.rdat2),
    .\rfif.rdat1 (rfif.rdat1),
    .\rfif.wdat (rfif.wdat),
    .\rfif.rsel2 (rfif.rsel2),
    .\rfif.rsel1 (rfif.rsel1),
    .\rfif.wsel (rfif.wsel),
    .\rfif.WEN (rfif.WEN),
    .\nRST (nRST),
    .\CLK (CLK)
  );
`endif

endmodule



program test(input logic CLK,
output logic nRST,
register_file_if.tb rfif);

parameter PERIOD = 10;

task reset_dut;
begin
  nRST = 0;
  @(posedge CLK);
  @(posedge CLK);
  @(negedge CLK);

  nRST = 1;
  @(posedge CLK);
  @(posedge CLK);

end
endtask


task write_reg;
input logic [4:0] reg_num;
input logic [31:0] reg_value;

begin
  rfif.wsel = reg_num;
  rfif.wdat = reg_value;
  @(negedge CLK);
end
endtask

task read_reg;
input logic [4:0] reg_num1;
input logic [4:0] reg_num2;

begin
  rfif.rsel1 = reg_num1;
  rfif.rsel2 = reg_num2;
  @(negedge CLK);
end
endtask

initial begin

  rfif.WEN = 0;
  rfif.wsel = 0;
  rfif.rsel1 = 0;
  rfif.rsel2 = 0;
  rfif.wdat = 0;
  nRST = 1;
  reset_dut;

  rfif.WEN = 1;

  rfif.rsel1 = 'd1;
  rfif.rsel2 = 'd2;
  @(negedge CLK);

  write_reg('d1, 'hAA);
  write_reg('d2, 'hBB);
  write_reg('d3, 'hCC);
  write_reg('d4, 'hDD);
  write_reg('d5, 'hEE);
  write_reg('d6, 'hFF);
  write_reg('d0, 'hEE);
  read_reg('d3,'d4);
  read_reg('d5,'d6);

  rfif.WEN = 0;
  write_reg('d1, 'hFF);
  read_reg('d1, 'd2);

  rfif.WEN = 1;
  write_reg('d1,'h22);
  write_reg('d0,'h50);
  

  $finish;

  end
endprogram
